module alu(inter.prakash face);
  always @(*) begin
  	face.out = face.a + face.b;
  end 
endmodule
